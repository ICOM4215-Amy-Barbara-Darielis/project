// Code your testbench here
// or browse Examples
/***
11100000100000100101000000000101
11100010010100110011000000000001
00011010111111111111111111111101
11100101110000010101000000000011
11011011000000000000000000000001
00000000000000000000000000000000
00000000000000000000000000000000
00000000000000000000000000000000
00000000000000000000000000000000**/

/*
1110000 0100 000100101000000000101 (ADD R5,R2,R5)
1110 001 0010 100110011000000000001 (SUBS R3,R3, #1)
0001101 0111 111111111111111111101 (BNE -3)

1110010 1110 000010101000000000011 (STRB R5, [R1,#3])

1101101 1000 000000000000000000001 (BLLE +2)
0000000 0000 000000000000000000000 (NOP)
*/
